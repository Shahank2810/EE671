VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO buffer
  CLASS BLOCK ;
  FOREIGN buffer ;
  ORIGIN 0.170 0.030 ;
  SIZE 4.580 BY 2.470 ;
  PIN Vss
    ANTENNADIFFAREA 0.604800 ;
    PORT
      LAYER li1 ;
        RECT 0.420 1.890 1.080 2.310 ;
        RECT 2.710 1.890 3.370 2.310 ;
      LAYER met1 ;
        RECT 0.420 2.280 0.840 2.310 ;
        RECT 2.710 2.280 3.130 2.310 ;
        RECT -0.170 1.950 4.410 2.280 ;
        RECT 0.420 1.890 0.840 1.950 ;
        RECT 2.710 1.890 3.130 1.950 ;
    END
  END Vss
  PIN Vdd
    ANTENNADIFFAREA 1.022000 ;
    PORT
      LAYER nwell ;
        RECT 0.260 0.400 4.060 1.500 ;
      LAYER li1 ;
        RECT 0.440 0.590 1.100 1.320 ;
        RECT 2.730 0.590 3.390 1.320 ;
      LAYER met1 ;
        RECT 0.440 1.060 0.840 1.320 ;
        RECT 2.730 1.060 3.130 1.320 ;
        RECT -0.170 0.730 4.410 1.060 ;
        RECT 0.440 0.590 0.840 0.730 ;
        RECT 2.730 0.590 3.130 0.730 ;
    END
  END Vdd
  PIN A
    ANTENNAGATEAREA 0.172500 ;
    PORT
      LAYER li1 ;
        RECT 1.000 0.240 1.320 0.310 ;
        RECT -0.170 0.000 1.320 0.240 ;
        RECT 1.000 -0.030 1.320 0.000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 0.345000 ;
    PORT
      LAYER li1 ;
        RECT 3.620 1.780 3.880 2.310 ;
        RECT 3.620 1.540 4.410 1.780 ;
        RECT 3.620 0.590 3.880 1.540 ;
        RECT 4.120 0.000 4.410 1.540 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 1.330 1.780 1.590 2.310 ;
        RECT 1.330 1.540 2.120 1.780 ;
        RECT 1.330 0.590 1.590 1.540 ;
        RECT 1.830 0.240 2.120 1.540 ;
        RECT 3.290 0.240 3.610 0.310 ;
        RECT 1.830 0.000 3.610 0.240 ;
        RECT 3.290 -0.030 3.610 0.000 ;
  END
END buffer
END LIBRARY

