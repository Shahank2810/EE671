magic
tech sky130A
timestamp 1725988179
<< nwell >>
rect 175 40 293 150
<< locali >>
rect -17 0 -1 24
rect 412 0 441 18
<< metal1 >>
rect -17 195 -2 228
rect -17 73 -2 106
use Inv  Inv_0 ~/shas
timestamp 1725987889
transform 1 0 115 0 1 172
box -132 -175 97 72
use Inv  Inv_1
timestamp 1725987889
transform 1 0 344 0 1 172
box -132 -175 97 72
<< labels >>
rlabel metal1 -17 211 -16 211 3 Vss
port 1 e
rlabel metal1 -17 88 -17 88 3 Vdd
port 2 e
rlabel locali -17 11 -17 11 3 A
port 3 e
rlabel locali 426 0 426 0 1 Y
port 4 n
<< end >>
