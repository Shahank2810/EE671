* NGSPICE file created from invx2.ext - technology: sky130A

.subckt invx2 Vdd Y A Vss
X0 Y A Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0.45 pd=3.6 as=0.45 ps=3.6 w=1.5 l=0.15
**devattr s=4500,360 d=4500,360
X1 Y A Vss Vss sky130_fd_pr__nfet_01v8 ad=0.252 pd=2.28 as=0.252 ps=2.28 w=0.84 l=0.15
**devattr s=2520,228 d=2520,228
.ends

